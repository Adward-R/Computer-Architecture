//Macro.vh
//macro definitions

//ALU CONTROL CODES
`define ALU_CTL_AND	3'b000
`define ALU_CTL_OR	3'b001
`define ALU_CTL_ADD	3'b010
`define ALU_CTL_SUB	3'b110
`define ALU_CTL_SLT	3'b111