`timescale 1ns / 1ps

`define DEBUG

// uncomment below macros when simulating this project
//`define SIMULATING